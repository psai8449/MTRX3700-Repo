//fsm

module fsm (
	input logic CLOCK,
	input logic [3:0] buttons
);




endmodule

