//motor_ctrl

module motor_ctrl 
(
	output logic [3:0] left,
	output logic [3:0] right,
	
	input logic [7:0] command
);

always_comb begin:

	case(command)
		

end


endmodule
