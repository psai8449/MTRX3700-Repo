//IR interpreter

// converts IR signals to commands the project will understand

module ir_interpreter (
	input logic [31:0] ir_input,
	
	output logic [7:0] ir_command
);



endmodule


